// File Name	: not_gate.v 
// Author		: Sibi Ravichandran
// Date			: 21-May-2020
// Description	: The function of this component is to perform NOT operation on a binary input.
//  Input-1 Output
//	  0		   1
//	  1		   0

// *********************************START OF CODE ********************************************************

module NOT (output Y, input A);
    not(Y, A); 
endmodule

// *********************************END OF CODE **********************************************************